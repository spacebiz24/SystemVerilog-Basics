class packet;
    randc bit [1:0]D;
    randc bit sel;
    bit rst;
    bit Q;
    
    // constraint random {D <= 3; sel <= 1;}
endclass
