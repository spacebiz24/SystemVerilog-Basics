class packet;
    rand bit [1:0]D;
    rand bit sel;
    bit rst;
    bit Q;
    
    // constraint random {D <= 3; sel <= 1;}
endclass
