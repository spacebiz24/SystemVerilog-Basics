`timescale 1ns / 1ps

interface DUT_interface();
  	logic [16]Operand1, Operand2;
  	logic [4]OpCode;
	logic [32]Result;
endinterface
